
module imem(input logic [5:0] a,
            output logic [18:0] rd);
  
  logic [18:0] IRAM [63:0];
  
  initial begin
    $readmemh("memfile1.hex",IRAM);
  end
  
  initial begin
//     IRAM[0]=19'b000_0011_1000_0100_0010;    // addi x2,x0,7
//     IRAM[1]=19'b000_0010_1000_0110_0010;    // addi x3,x0,5
//     IRAM[2]=19'b000_1101_0011_1000_0001;    // mul x4,x3,x2   // checked
    
//     IRAM[0]=19'b000_0011_1000_0100_0010;    // addi x2,x0,7
//     IRAM[1]=19'b000_0010_1000_0110_0010;    // addi x3,x0,5
//     IRAM[2]=19'b010_1101_1010_1010_0001;    // rem x5,x2,x3
//     IRAM[3]=19'b001_0001_1010_1100_0001;    // div x6,x2,x3
//     IRAM[4]=19'b000_1001_1010_1110_0001;    // sub x7,x2,x3    // checked
    
//     IRAM[0]=19'b000_0011_1000_0100_0010;    // addi x2,x0,7
//     IRAM[1]=19'b000_0010_1000_0110_0010;    // addi x3,x0,5
//     IRAM[2]=19'b001_0100_0010_0100_0001;    // inc x2
//     IRAM[3]=19'b001_1000_0011_0110_0001;    // dec x3          // checked
    
//     IRAM[0]=19'b000_0011_1000_0100_0010;    // addi x2,x0,7
//     IRAM[1]=19'b000_0010_1000_0110_0010;    // addi x3,x0,5
//     IRAM[2]=19'b001_1101_1010_1010_0001;    // and x5,x2,x3
//     IRAM[3]=19'b010_0001_1010_1000_0001;    // or x4,x2,x3
//     IRAM[4]=19'b010_0101_1010_1100_0001;    // xor x6,x2,x3
//     IRAM[5]=19'b010_1000_0110_1100_0001;    // not x6          // checked
    
//     IRAM[0]=19'b000_0011_1000_0100_0010;    // addi x2,x0,7
//     IRAM[1]=19'b000_0001_0000_0110_0010;    // addi x3,x0,2
//     IRAM[2]=19'b011_0001_1010_1010_0001;    // slt x5,x2,x3
//     IRAM[3]=19'b011_0101_1010_1100_0001;    // sll x6,x2,x3
//     IRAM[4]=19'b011_1001_1010_1110_0001;    // srl x7,x2,x3
//     IRAM[5]=19'b011_1101_1010_1000_0001;    // sra x4,x2,x3     // checked
    
//     IRAM[0]=19'b000_0100_1000_0010_0010;    // addi x1,x0,9
//     IRAM[1]=19'b000_0010_1001_0100_0110;    // muli x2,x1,5
//     IRAM[2]=19'b000_0101_0001_0110_1010;    // andi x3,x1,a
//     IRAM[3]=19'b000_0001_1001_1010_0111;    // divi x5,x1,3     // checked
    
//     IRAM[0]=19'b000_0010_0000_0110_0010;    // addi x3,x0,4
//     IRAM[1]=19'b010_0001_1000_1000_0100;    // sw x3,68(x0)
//     IRAM[2]=19'b010_0010_0000_0100_0011;    // lw x2,68(x0)     // checked
    
//     IRAM[0]=19'b000_0100_1000_0110_0010;    //       addi x3,x0,9
//     IRAM[1]=19'b000_0100_1000_1000_0010;    //       addi x4,x0,9
//     IRAM[2]=19'b000_0010_0011_1100_1000;    //       beq x3,x4,done
//     IRAM[3]=19'b000_0010_1011_1010_1010;    //       andi x5,x3,5
//     IRAM[4]=19'b000_0010_0011_1000_1000;    //       add x1,x3,x4
//     IRAM[5]=19'b000_0101_0011_1110_0110;   // done: muli x7,x3,a// checked
    
//     IRAM[0]=19'b000_0010_1000_0100_0010; //        addi x1,x0,5
//     IRAM[1]=19'b000_0000_1001_0101_0000; //        jal x2,target
//     IRAM[2]=19'b000_0100_1000_0110_0010; //        addi x3,x0,9
//     IRAM[3]=19'b000_0001_1000_1010_0010; //target: addi x5,x0,3 // checked
    
//     IRAM[0]=19'b000_0100_1000_0110_0010;    //       addi x3,x0,9
//     IRAM[1]=19'b000_0010_1000_1000_0010;    //       addi x4,x0,5
//     IRAM[2]=19'b000_0010_0011_1100_1110;    //       bne x3,x4,done
//     IRAM[3]=19'b000_0010_1011_1010_1010;    //       andi x5,x3,5
//     IRAM[4]=19'b000_0010_0011_1000_1000;    //       add x1,x3,x4
//     IRAM[5]=19'b000_0101_0011_1110_0110;   // done: muli x7,x3,a// checked
  end
  
  assign rd = IRAM[a];
endmodule